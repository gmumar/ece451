magic
tech scmos
use /nfs/ug/homes-0/s/syedazaa/ECE451/git_folder/ece451/lab2/OneBit_Slice.lvs /nfs/ug/homes-0/s/syedazaa/ECE451/git_folder/ece451/lab2/OneBit_Slice.lvs_0
transform 1 0 0 0 1 0
box 0 0 10 10
<< error_s >>
rect 963 645 966 648
<< labels >>
rlabel space 963 645 963 645 2 [S]gnd
<< error_s >>
rect 436 760 439 763
<< labels >>
rlabel space 436 760 436 760 2 [S]gnd
<< error_s >>
rect 417 760 420 763
<< labels >>
rlabel space 417 760 417 760 2 [S]gnd
<< error_s >>
rect 377 760 380 763
<< labels >>
rlabel space 377 760 377 760 2 [S]gnd
<< error_s >>
rect 357 760 360 763
<< labels >>
rlabel space 357 760 357 760 2 [S]gnd
<< error_s >>
rect -363 766 -360 769
<< labels >>
rlabel space -363 766 -363 766 2 [S]gnd
<< error_s >>
rect -442 766 -439 769
<< labels >>
rlabel space -442 766 -442 766 2 [S]gnd
<< error_s >>
rect -462 766 -459 769
<< labels >>
rlabel space -462 766 -462 766 2 [S]gnd
<< error_s >>
rect -573 772 -570 775
<< labels >>
rlabel space -573 772 -573 772 2 [S]gnd
<< error_s >>
rect -736 766 -733 769
<< labels >>
rlabel space -736 766 -736 766 2 [S]gnd
<< error_s >>
rect -815 766 -812 769
<< labels >>
rlabel space -815 766 -815 766 2 [S]gnd
<< error_s >>
rect -835 766 -832 769
<< labels >>
rlabel space -835 766 -835 766 2 [S]gnd
<< error_s >>
rect -1132 762 -1129 765
<< labels >>
rlabel space -1132 762 -1132 762 2 [S]gnd
<< error_s >>
rect -1448 762 -1445 765
<< labels >>
rlabel space -1448 762 -1448 762 2 [S]gnd
<< error_s >>
rect -1764 762 -1761 765
<< labels >>
rlabel space -1764 762 -1764 762 2 [S]gnd
<< error_s >>
rect -2079 762 -2076 765
<< labels >>
rlabel space -2079 762 -2079 762 2 [S]gnd
<< error_s >>
rect -1448 782 -1445 785
<< labels >>
rlabel space -1448 782 -1448 782 2 [S]gnd
<< error_s >>
rect -1764 782 -1761 785
<< labels >>
rlabel space -1764 782 -1764 782 2 [S]gnd
<< error_s >>
rect -2079 782 -2076 785
<< labels >>
rlabel space -2079 782 -2079 782 2 [S]gnd
<< error_s >>
rect -1448 762 -1445 765
<< labels >>
rlabel space -1448 762 -1448 762 4 [G]RegFile_79/RamCell_4/#fet_75/d
<< error_s >>
rect -1448 782 -1445 785
<< labels >>
rlabel space -1448 782 -1448 782 2 [S]RegFile_79/RamCell_4/#fet_75/d
<< error_s >>
rect -1516 762 -1513 765
<< labels >>
rlabel space -1516 762 -1516 762 4 [G]RegFile_79/RamCell_4/#fet_75/d
<< error_s >>
rect -1516 782 -1513 785
<< labels >>
rlabel space -1516 782 -1516 782 2 [S]RegFile_79/RamCell_4/#fet_75/d
<< error_s >>
rect -2202 749 -2199 752
<< labels >>
rlabel space -2202 749 -2202 749 2 [S]RegFile_79/RamCell_45/#fet!-type!pfet!-width!2.0_0/s
<< error_s >>
rect -2202 769 -2199 772
<< labels >>
rlabel space -2202 769 -2202 769 2 [S]RegFile_79/RamCell_45/#fet!-type!pfet!-width!2.0_0/s
<< error_s >>
rect -2079 782 -2076 785
<< labels >>
rlabel space -2079 782 -2079 782 4 [G]RegFile_79/RamCell_45/#fet!-type!pfet!-width!2.0_0/s
<< error_s >>
rect -2147 743 -2144 746
<< labels >>
rlabel space -2147 743 -2147 743 2 [S]RegFile_79/RamCell_45/#fet!-type!pfet!-width!2.0_0/s
<< error_s >>
rect -2147 782 -2144 785
<< labels >>
rlabel space -2147 782 -2147 782 4 [G]RegFile_79/RamCell_45/#fet!-type!pfet!-width!2.0_0/s
<< error_s >>
rect -1570 749 -1567 752
<< labels >>
rlabel space -1570 749 -1570 749 2 [S]RegFile_79/RamCell_4/#fet!-type!pfet!-width!2.0_0/s
<< error_s >>
rect -1570 769 -1567 772
<< labels >>
rlabel space -1570 769 -1570 769 2 [S]RegFile_79/RamCell_4/#fet!-type!pfet!-width!2.0_0/s
<< error_s >>
rect -1448 782 -1445 785
<< labels >>
rlabel space -1448 782 -1448 782 4 [G]RegFile_79/RamCell_4/#fet!-type!pfet!-width!2.0_0/s
<< error_s >>
rect -1516 743 -1513 746
<< labels >>
rlabel space -1516 743 -1516 743 2 [S]RegFile_79/RamCell_4/#fet!-type!pfet!-width!2.0_0/s
<< error_s >>
rect -1516 782 -1513 785
<< labels >>
rlabel space -1516 782 -1516 782 4 [G]RegFile_79/RamCell_4/#fet!-type!pfet!-width!2.0_0/s
<< error_s >>
rect -1516 743 -1513 746
<< labels >>
rlabel space -1516 743 -1516 743 4 [G]notFBEn[2]
<< error_s >>
rect -1764 762 -1761 765
<< labels >>
rlabel space -1764 762 -1764 762 2 [S]RegFile_79/RamCell_2/#fet_87/s
<< error_s >>
rect -1886 769 -1883 772
<< labels >>
rlabel space -1886 769 -1886 769 2 [S]RegFile_79/RamCell_2/#fet_87/s
<< error_s >>
rect -1885 810 -1882 813
<< labels >>
rlabel space -1885 810 -1885 810 2 [S]RegFile_79/RamCell_2/#fet_87/s
<< error_s >>
rect -1885 829 -1882 832
<< labels >>
rlabel space -1885 829 -1885 829 2 [S]RegFile_79/RamCell_2/#fet_87/s
<< error_s >>
rect -1831 743 -1828 746
<< labels >>
rlabel space -1831 743 -1831 743 2 [S]RegFile_79/RamCell_2/#fet_87/s
<< error_s >>
rect -1831 762 -1828 765
<< labels >>
rlabel space -1831 762 -1831 762 2 [S]RegFile_79/RamCell_2/#fet_87/s
<< error_s >>
rect -1448 762 -1445 765
<< labels >>
rlabel space -1448 762 -1448 762 2 [S]RegFile_79/RamCell_4/#fet_87/s
<< error_s >>
rect -1570 769 -1567 772
<< labels >>
rlabel space -1570 769 -1570 769 2 [S]RegFile_79/RamCell_4/#fet_87/s
<< error_s >>
rect -1570 810 -1567 813
<< labels >>
rlabel space -1570 810 -1570 810 2 [S]RegFile_79/RamCell_4/#fet_87/s
<< error_s >>
rect -1570 829 -1567 832
<< labels >>
rlabel space -1570 829 -1570 829 2 [S]RegFile_79/RamCell_4/#fet_87/s
<< error_s >>
rect -1516 743 -1513 746
<< labels >>
rlabel space -1516 743 -1516 743 2 [S]RegFile_79/RamCell_4/#fet_87/s
<< error_s >>
rect -1516 762 -1513 765
<< labels >>
rlabel space -1516 762 -1516 762 2 [S]RegFile_79/RamCell_4/#fet_87/s
<< error_s >>
rect 963 690 966 693
<< labels >>
rlabel space 963 690 963 690 2 [S]vdd
<< error_s >>
rect -1200 762 -1197 765
<< labels >>
rlabel space -1200 762 -1200 762 2 [S]vdd
<< error_s >>
rect -1516 762 -1513 765
<< labels >>
rlabel space -1516 762 -1516 762 2 [S]vdd
<< error_s >>
rect -1831 762 -1828 765
<< labels >>
rlabel space -1831 762 -1831 762 2 [S]vdd
<< error_s >>
rect -2147 762 -2144 765
<< labels >>
rlabel space -2147 762 -2147 762 2 [S]vdd
<< error_s >>
rect -1516 782 -1513 785
<< labels >>
rlabel space -1516 782 -1516 782 2 [S]vdd
<< error_s >>
rect -1831 782 -1828 785
<< labels >>
rlabel space -1831 782 -1831 782 2 [S]vdd
<< error_s >>
rect -2147 782 -2144 785
<< labels >>
rlabel space -2147 782 -2147 782 2 [S]vdd
<< error_s >>
rect 417 812 420 815
<< labels >>
rlabel space 417 812 417 812 2 [S]vdd
<< error_s >>
rect 377 812 380 815
<< labels >>
rlabel space 377 812 377 812 2 [S]vdd
<< error_s >>
rect 357 812 360 815
<< labels >>
rlabel space 357 812 357 812 2 [S]vdd
<< error_s >>
rect -570 827 -567 830
<< labels >>
rlabel space -570 827 -570 827 2 [S]vdd
<< error_s >>
rect -943 827 -940 830
<< labels >>
rlabel space -943 827 -943 827 2 [S]vdd
<< error_s >>
rect 418 882 421 885
<< labels >>
rlabel space 418 882 418 882 2 [S]vdd
<< error_s >>
rect 377 882 380 885
<< labels >>
rlabel space 377 882 377 882 2 [S]vdd
<< error_s >>
rect 357 882 360 885
<< labels >>
rlabel space 357 882 357 882 2 [S]vdd
<< error_s >>
rect -363 855 -360 858
<< labels >>
rlabel space -363 855 -363 855 2 [S]vdd
<< error_s >>
rect -442 855 -439 858
<< labels >>
rlabel space -442 855 -442 855 2 [S]vdd
<< error_s >>
rect -462 855 -459 858
<< labels >>
rlabel space -462 855 -462 855 2 [S]vdd
<< error_s >>
rect -736 855 -733 858
<< labels >>
rlabel space -736 855 -736 855 2 [S]vdd
<< error_s >>
rect -815 855 -812 858
<< labels >>
rlabel space -815 855 -815 855 2 [S]vdd
<< error_s >>
rect -835 855 -832 858
<< labels >>
rlabel space -835 855 -835 855 2 [S]vdd
<< error_s >>
rect -2373 852 -2370 855
<< labels >>
rlabel space -2373 852 -2373 852 2 [S]vdd
<< error_s >>
rect -2393 852 -2390 855
<< labels >>
rlabel space -2393 852 -2393 852 2 [S]vdd
<< error_s >>
rect -892 752 -889 755
<< labels >>
rlabel space -892 752 -892 752 2 [S]D
<< error_s >>
rect -1254 749 -1251 752
<< labels >>
rlabel space -1254 749 -1254 749 2 [S]D
<< error_s >>
rect -1254 749 -1251 752
<< labels >>
rlabel space -1254 749 -1254 749 2 [S]D
<< error_s >>
rect -1570 749 -1567 752
<< labels >>
rlabel space -1570 749 -1570 749 2 [S]D
<< error_s >>
rect -1886 749 -1883 752
<< labels >>
rlabel space -1886 749 -1886 749 2 [S]D
<< error_s >>
rect -2202 749 -2199 752
<< labels >>
rlabel space -2202 749 -2202 749 2 [S]D
<< error_s >>
rect -1132 762 -1129 765
<< labels >>
rlabel space -1132 762 -1132 762 2 [S]D
<< error_s >>
rect -1132 762 -1129 765
<< labels >>
rlabel space -1132 762 -1132 762 2 [S]D
<< error_s >>
rect -946 772 -943 775
<< labels >>
rlabel space -946 772 -946 772 2 [S]D
<< error_s >>
rect -1254 769 -1251 772
<< labels >>
rlabel space -1254 769 -1254 769 2 [S]D
<< error_s >>
rect -1254 769 -1251 772
<< labels >>
rlabel space -1254 769 -1254 769 2 [S]D
<< error_s >>
rect -2533 785 -2530 788
<< labels >>
rlabel space -2533 785 -2533 785 2 [S]D
<< error_s >>
rect -1254 810 -1251 813
<< labels >>
rlabel space -1254 810 -1254 810 2 [S]D
<< error_s >>
rect -1254 810 -1251 813
<< labels >>
rlabel space -1254 810 -1254 810 2 [S]D
<< error_s >>
rect -1570 810 -1567 813
<< labels >>
rlabel space -1570 810 -1570 810 2 [S]D
<< error_s >>
rect -1885 810 -1882 813
<< labels >>
rlabel space -1885 810 -1885 810 2 [S]D
<< error_s >>
rect -2201 810 -2198 813
<< labels >>
rlabel space -2201 810 -2201 810 2 [S]D
<< error_s >>
rect -1254 829 -1251 832
<< labels >>
rlabel space -1254 829 -1254 829 2 [S]D
<< error_s >>
rect -2537 852 -2534 855
<< labels >>
rlabel space -2537 852 -2537 852 2 [S]D
<< error_s >>
rect -1200 743 -1197 746
<< labels >>
rlabel space -1200 743 -1200 743 2 [S]D
<< error_s >>
rect -1200 743 -1197 746
<< labels >>
rlabel space -1200 743 -1200 743 2 [S]D
<< error_s >>
rect -1200 743 -1197 746
<< labels >>
rlabel space -1200 743 -1200 743 2 [S]D
<< error_s >>
rect -1200 762 -1197 765
<< labels >>
rlabel space -1200 762 -1200 762 2 [S]D
<< error_s >>
rect -1200 762 -1197 765
<< labels >>
rlabel space -1200 762 -1200 762 2 [S]D
<< error_s >>
rect -2617 785 -2614 788
<< labels >>
rlabel space -2617 785 -2617 785 2 [S]D
<< error_s >>
rect -2373 852 -2370 855
<< labels >>
rlabel space -2373 852 -2373 852 2 [S]D
<< error_s >>
rect -2617 852 -2614 855
<< labels >>
rlabel space -2617 852 -2617 852 2 [S]D
<< error_s >>
rect -1200 762 -1197 765
<< labels >>
rlabel space -1200 762 -1200 762 8 D:
<< error_s >>
rect -1516 743 -1513 746
<< labels >>
rlabel space -1516 743 -1516 743 8 D:
<< error_s >>
rect -1516 762 -1513 765
<< labels >>
rlabel space -1516 762 -1516 762 8 D:
<< error_s >>
rect -1516 782 -1513 785
<< labels >>
rlabel space -1516 782 -1516 782 8 D:
<< error_s >>
rect -1200 743 -1197 746
<< labels >>
rlabel space -1200 743 -1200 743 8 D:
<< error_s >>
rect -1448 782 -1445 785
<< labels >>
rlabel space -1448 782 -1448 782 8 D:
<< error_s >>
rect -1448 762 -1445 765
<< labels >>
rlabel space -1448 762 -1448 762 8 D:
<< error_s >>
rect -1132 762 -1129 765
<< labels >>
rlabel space -1132 762 -1132 762 8 D:
<< end >>
