magic
tech scmos
use /nfs/ug/homes-2/u/umarghul/ece451/lab2/RamCell.lvs /nfs/ug/homes-2/u/umarghul/ece451/lab2/RamCell.lvs_0
transform 1 0 0 0 1 0
box 0 0 10 10
<< end >>
