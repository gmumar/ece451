* FILE: test_inv.sp

********************** begin header *****************************

* Sample Header file for Generic 2.5V 0.25 um process (g25)

.OPTIONS post ACCT OPTS lvltim=2
.OPTIONS post_version=9007

**################################################
* Only Typical/Typical models included
* NEED TO CHANGE ${MMI_TOOLS} TO BE PHYSICAL PATH
.include '/cad2/mmi_local/sue/g25.mod'
* NOTE: these are contrived spice models
**################################################

.param  arean(w,sdd) = '(w*sdd*1p)'
.param  areap(w,sdd) = '(w*sdd*1p)'
* Setup either one or the other of the following
* For ACM=0,2,10,12 fet models
.param  perin(w,sdd) = '(2u*(w+sdd))'
.param  perip(w,sdd) = '(2u*(w+sdd))'
* For ACM=3,13 fet models
*.param  perin(w,sdd) = '(1u*(w+2*sdd))'
*.param  perip(w,sdd) = '(1u*(w+2*sdd))'

.param ln_min   =  0.25u
.param lp_min   =  0.25u

* used in source/drain area/perimeter calculation
.param sdd        =  0.95

.PARAM vddp=2.5		$ VDD voltage

VDD vdd 0 DC vddp 

.TEMP 105
.TRAN 10p 16n
*********************** end header ******************************

* SPICE netlist for "test_inv" generated by MMI_SUE5.5.4 on Mon Jan 12 
*+ 11:18:12 AM EST 2015.

.SUBCKT Counter OUT1 OUT2 
V_1 OUT2 GND pulse 0 vddp 0ns 200ps 200ps 3ns 6ns 
V_2 OUT1 GND pulse 0 vddp 0ns 200ps 200ps 6ns 12ns 
.ENDS	$ Counter

.SUBCKT inv A out 
M_1 out A vdd vdd p W='2*1u' L=lp_min ad='areap(2,sdd)' 
+ as='areap(2,sdd)' pd='perip(2,sdd)' ps='perip(2,sdd)' 
M_2 out A gnd gnd n W='1*1u' L=ln_min ad='arean(1,sdd)' 
+ as='arean(1,sdd)' pd='perin(1,sdd)' ps='perin(1,sdd)' 
.ENDS	$ inv

* start main CELL test_inv
* .SUBCKT test_inv  
XCounter net_1 uc_net_2 Counter 
Xinv net_1 uc_net_3 inv 
* .ENDS	$ test_inv

.GLOBAL gnd vdd

.END

