magic
tech scmos
use /nfs/ug/homes-2/u/umarghul/ece451/lab2/ALU.lvs /nfs/ug/homes-2/u/umarghul/ece451/lab2/ALU.lvs_0
transform 1 0 0 0 1 0
box 0 0 10 10
<< error_s >>
rect -975 224 -972 227
<< labels >>
rlabel space -975 224 -975 224 2 [S]Func_82/Y
<< error_s >>
rect -975 244 -972 247
<< labels >>
rlabel space -975 244 -975 244 2 [S]Func_82/Y
<< error_s >>
rect -975 313 -972 316
<< labels >>
rlabel space -975 313 -975 313 2 [S]Func_82/Y
<< error_s >>
rect -975 332 -972 335
<< labels >>
rlabel space -975 332 -975 332 2 [S]Func_82/Y
<< error_s >>
rect -326 236 -323 239
<< labels >>
rlabel space -326 236 -326 236 2 [S]Carry_99/notCi
<< error_s >>
rect -346 236 -343 239
<< labels >>
rlabel space -346 236 -346 236 2 [S]Carry_99/notCi
<< error_s >>
rect -364 358 -361 361
<< labels >>
rlabel space -364 358 -364 358 2 [S]Carry_99/notCi
<< error_s >>
rect 43 224 46 227
<< labels >>
rlabel space 43 224 43 224 2 [S]TFunc_95/Y
<< error_s >>
rect 43 244 46 247
<< labels >>
rlabel space 43 244 43 244 2 [S]TFunc_95/Y
<< error_s >>
rect 43 312 46 315
<< labels >>
rlabel space 43 312 43 312 2 [S]TFunc_95/Y
<< error_s >>
rect 43 332 46 335
<< labels >>
rlabel space 43 332 43 332 2 [S]TFunc_95/Y
<< error_s >>
rect -220 224 -217 227
<< labels >>
rlabel space -220 224 -220 224 2 [S]TFunc_95/Y
<< error_s >>
rect -220 244 -217 247
<< labels >>
rlabel space -220 244 -220 244 2 [S]TFunc_95/Y
<< error_s >>
rect -220 312 -217 315
<< labels >>
rlabel space -220 312 -220 312 2 [S]TFunc_95/Y
<< error_s >>
rect -220 332 -217 335
<< labels >>
rlabel space -220 332 -220 332 2 [S]TFunc_95/Y
<< error_s >>
rect -346 236 -343 239
<< labels >>
rlabel space -346 236 -346 236 2 [S]gnd
<< error_s >>
rect -366 236 -363 239
<< labels >>
rlabel space -366 236 -366 236 2 [S]gnd
<< error_s >>
rect -406 236 -403 239
<< labels >>
rlabel space -406 236 -406 236 2 [S]gnd
<< error_s >>
rect -425 236 -422 239
<< labels >>
rlabel space -425 236 -425 236 2 [S]gnd
<< error_s >>
rect 43 298 46 301
<< labels >>
rlabel space 43 298 43 298 4 [G]TFunc_95/notR
<< error_s >>
rect 43 332 46 335
<< labels >>
rlabel space 43 332 43 332 4 [G]TFunc_95/notR
<< error_s >>
rect -220 224 -217 227
<< labels >>
rlabel space -220 224 -220 224 4 [G]TFunc_95/notR
<< error_s >>
rect -220 258 -217 261
<< labels >>
rlabel space -220 258 -220 258 4 [G]TFunc_95/notR
<< error_s >>
rect 43 209 46 212
<< labels >>
rlabel space 43 209 43 209 2 [S]TFunc_95/X[3]
<< error_s >>
rect -220 209 -217 212
<< labels >>
rlabel space -220 209 -220 209 2 [S]TFunc_95/X[3]
<< error_s >>
rect 43 347 46 350
<< labels >>
rlabel space 43 347 43 347 2 [S]TFunc_95/X[0]
<< error_s >>
rect -220 347 -217 350
<< labels >>
rlabel space -220 347 -220 347 2 [S]TFunc_95/X[0]
<< error_s >>
rect -366 288 -363 291
<< labels >>
rlabel space -366 288 -366 288 2 [S]vdd
<< error_s >>
rect -406 288 -403 291
<< labels >>
rlabel space -406 288 -406 288 2 [S]vdd
<< error_s >>
rect -425 288 -422 291
<< labels >>
rlabel space -425 288 -425 288 2 [S]vdd
<< error_s >>
rect -364 358 -361 361
<< labels >>
rlabel space -364 358 -364 358 2 [S]vdd
<< error_s >>
rect -405 358 -402 361
<< labels >>
rlabel space -405 358 -405 358 2 [S]vdd
<< error_s >>
rect -425 358 -422 361
<< labels >>
rlabel space -425 358 -425 358 2 [S]vdd
<< error_s >>
rect -366 236 -363 239
<< labels >>
rlabel space -366 236 -366 236 4 [G]Carry_99/#fet_83/d
<< error_s >>
rect -366 288 -363 291
<< labels >>
rlabel space -366 288 -366 288 4 [G]Carry_99/#fet_83/d
<< error_s >>
rect -405 358 -402 361
<< labels >>
rlabel space -405 358 -405 358 2 [S]Carry_99/#fet_83/d
<< error_s >>
rect 43 258 46 261
<< labels >>
rlabel space 43 258 43 258 4 [G]TFunc_95/notS
<< error_s >>
rect 43 347 46 350
<< labels >>
rlabel space 43 347 43 347 4 [G]TFunc_95/notS
<< error_s >>
rect -220 209 -217 212
<< labels >>
rlabel space -220 209 -220 209 4 [G]TFunc_95/notS
<< error_s >>
rect -220 298 -217 301
<< labels >>
rlabel space -220 298 -220 298 4 [G]TFunc_95/notS
<< end >>
